
library ieee;
use ieee.std_logic_1164.all;

entity sin_entity is
port ( address : in std_logic_vector(6 downto 0);
     data : out real );
end entity sin_entity;

architecture sin_arch of sin_entity is
type mem is array ( 0 to 99) of real;
constant my_rom : mem := (
0 =>0.0,
1 =>0.0627905195293134,
2 =>0.125333233564304,
3 =>0.187381314585725,
4 =>0.248689887164855,
5 =>0.309016994374947,
6 =>0.368124552684678,
7 =>0.425779291565073,
8 =>0.481753674101715,
9 =>0.535826794978997,
10 =>0.587785252292473,
11 =>0.637423989748690,
12 =>0.684547105928689,
13 =>0.728968627421412,
14 =>0.770513242775789,
15 =>0.809016994374948,
16 =>0.844327925502015,
17 =>0.876306680043864,
18 =>0.904827052466020,
19 =>0.929776485888251,
20 =>0.951056516295154,
21 =>0.968583161128631,
22 =>0.982287250728689,
23 =>0.992114701314478,
24 =>0.998026728428272,
25 =>1.0,
26 =>0.998026728428272,
27 =>0.992114701314478,
28 =>0.982287250728689,
29 =>0.968583161128631,
30 =>0.951056516295154,
31 =>0.929776485888252,
32 =>0.904827052466020,
33 =>0.876306680043864,
34 =>0.844327925502015,
35 =>0.809016994374948,
36 =>0.770513242775789,
37 =>0.728968627421411,
38 =>0.684547105928689,
39 =>0.637423989748690,
40 =>0.587785252292473,
41 =>0.535826794978997,
42 =>0.481753674101716,
43 =>0.425779291565073,
44 =>0.368124552684678,
45 =>0.309016994374948,
46 =>0.248689887164855,
47 =>0.187381314585725,
48 =>0.125333233564304,
49 =>0.0627905195293131,
50 =>1.01064309961486e-15,
51 =>-0.0627905195293125,
52 =>-0.125333233564303,
53 =>-0.187381314585724,
54 =>-0.248689887164854,
55 =>-0.309016994374946,
56 =>-0.368124552684678,
57 =>-0.425779291565072,
58 =>-0.481753674101715,
59 =>-0.535826794978996,
60 =>-0.587785252292473,
61 =>-0.637423989748689,
62 =>-0.684547105928688,
63 =>-0.728968627421411,
64 =>-0.770513242775789,
65 =>-0.809016994374947,
66 =>-0.844327925502015,
67 =>-0.876306680043864,
68 =>-0.904827052466019,
69 =>-0.929776485888251,
70 =>-0.951056516295154,
71 =>-0.968583161128631,
72 =>-0.982287250728689,
73 =>-0.992114701314478,
74 =>-0.998026728428272,
75 =>-1.0,
76 =>-0.998026728428272,
77 =>-0.992114701314478,
78 =>-0.982287250728689,
79 =>-0.968583161128631,
80 =>-0.951056516295154,
81 =>-0.929776485888252,
82 =>-0.904827052466020,
83 =>-0.876306680043864,
84 =>-0.844327925502016,
85 =>-0.809016994374948,
86 =>-0.770513242775790,
87 =>-0.728968627421412,
88 =>-0.684547105928689,
89 =>-0.637423989748690,
90 =>-0.587785252292474,
91 =>-0.535826794978997,
92 =>-0.481753674101715,
93 =>-0.425779291565074,
94 =>-0.368124552684679,
95 =>-0.309016994374948,
96 =>-0.248689887164855,
97 =>-0.187381314585726,
98 =>-0.125333233564305,
99 =>-0.0627905195293142);

begin
process (address)
begin
 case address is
 when "0000000" => data <= my_rom(0);
when "0000001" => data <= my_rom(1);
when "0000010" => data <= my_rom(2);
when "0000011" => data <= my_rom(3);
when "0000100" => data <= my_rom(4);
when "0000101" => data <= my_rom(5);
when "0000110" => data <= my_rom(6);
when "0000111" => data <= my_rom(7);
when "0001000" => data <= my_rom(8);
when "0001001" => data <= my_rom(9);
when "0001010" => data <= my_rom(10);
when "0001011" => data <= my_rom(11);
when "0001100" => data <= my_rom(12);
when "0001101" => data <= my_rom(13);
when "0001110" => data <= my_rom(14);
when "0001111" => data <= my_rom(15);
when "0010000" => data <= my_rom(16);
when "0010001" => data <= my_rom(17);
when "0010010" => data <= my_rom(18);
when "0010011" => data <= my_rom(19);
when "0010100" => data <= my_rom(20);
when "0010101" => data <= my_rom(21);
when "0010110" => data <= my_rom(22);
when "0010111" => data <= my_rom(23);
when "0011000" => data <= my_rom(24);
when "0011001" => data <= my_rom(25);
when "0011010" => data <= my_rom(26);
when "0011011" => data <= my_rom(27);
when "0011100" => data <= my_rom(28);
when "0011101" => data <= my_rom(29);
when "0011110" => data <= my_rom(30);
when "0011111" => data <= my_rom(31);
when "0100000" => data <= my_rom(32);
when "0100001" => data <= my_rom(33);
when "0100010" => data <= my_rom(34);
when "0100011" => data <= my_rom(35);
when "0100100" => data <= my_rom(36);
when "0100101" => data <= my_rom(37);
when "0100110" => data <= my_rom(38);
when "0100111" => data <= my_rom(39);
when "0101000" => data <= my_rom(40);
when "0101001" => data <= my_rom(41);
when "0101010" => data <= my_rom(42);
when "0101011" => data <= my_rom(43);
when "0101100" => data <= my_rom(44);
when "0101101" => data <= my_rom(45);
when "0101110" => data <= my_rom(46);
when "0101111" => data <= my_rom(47);
when "0110000" => data <= my_rom(48);
when "0110001" => data <= my_rom(49);
when "0110010" => data <= my_rom(50);
when "0110011" => data <= my_rom(51);
when "0110100" => data <= my_rom(52);
when "0110101" => data <= my_rom(53);
when "0110110" => data <= my_rom(54);
when "0110111" => data <= my_rom(55);
when "0111000" => data <= my_rom(56);
when "0111001" => data <= my_rom(57);
when "0111010" => data <= my_rom(58);
when "0111011" => data <= my_rom(59);
when "0111100" => data <= my_rom(60);
when "0111101" => data <= my_rom(61);
when "0111110" => data <= my_rom(62);
when "0111111" => data <= my_rom(63);
when "1000000" => data <= my_rom(64);
when "1000001" => data <= my_rom(65);
when "1000010" => data <= my_rom(66);
when "1000011" => data <= my_rom(67);
when "1000100" => data <= my_rom(68);
when "1000101" => data <= my_rom(69);
when "1000110" => data <= my_rom(70);
when "1000111" => data <= my_rom(71);
when "1001000" => data <= my_rom(72);
when "1001001" => data <= my_rom(73);
when "1001010" => data <= my_rom(74);
when "1001011" => data <= my_rom(75);
when "1001100" => data <= my_rom(76);
when "1001101" => data <= my_rom(77);
when "1001110" => data <= my_rom(78);
when "1001111" => data <= my_rom(79);
when "1010000" => data <= my_rom(80);
when "1010001" => data <= my_rom(81);
when "1010010" => data <= my_rom(82);
when "1010011" => data <= my_rom(83);
when "1010100" => data <= my_rom(84);
when "1010101" => data <= my_rom(85);
when "1010110" => data <= my_rom(86);
when "1010111" => data <= my_rom(87);
when "1011000" => data <= my_rom(88);
when "1011001" => data <= my_rom(89);
when "1011010" => data <= my_rom(90);
when "1011011" => data <= my_rom(91);
when "1011100" => data <= my_rom(92);
when "1011101" => data <= my_rom(93);
when "1011110" => data <= my_rom(94);
when "1011111" => data <= my_rom(95);
when "1100000" => data <= my_rom(96);
when "1100001" => data <= my_rom(97);
when "1100010" => data <= my_rom(98);
when "1100011" => data <= my_rom(99);

       when others => data <= 0.0;
         end case;
  end process;
end sin_arch;
