library ieee;
use ieee.std_logic_1164.all;

entity clocked_fsm is
	port(
		clk,reset : in std_logic;
		start: in std_logic; -- start waveform generation
		full: in std_logic; --Counter is Full
		P: out std_logic; --Counter Toggle?
		CC: out std_logic; -- Clear Clock
		CS: out std_logic;
		E: out std_logic;
		LP: out std_logic
	);
end entity clocked_fsm;

architecture clocked_fsm_arch of clocked_fsm is
	type waveform_state_type is (s0, s1, s2, s3);
	signal state_reg, state_next: waveform_state_type;
begin
	--State Register Logic
	process(clk, reset)
	begin
		-- Active Low FSM Reset?
		if (reset = '0') 
			then state_reg <=s0;
		elsif (clk'event and clk ='1') 
			then state_reg <= state_next;
		end if; 
	end process;

	--Next State Logic 
	process(state_reg, start)
	begin
		case state_reg is 
			when s0 => 
				if (start ='1') then state_next <= s1;
				else then state_next <= s0; end if;
			when s1 => 
				state_next <= s2;
			when s2 => 
				state_next <= s3;
			when s3 => 
				state_next <= s1;
		end case;
	end process;

	--Moore Output Logic
	process(state_reg)
	begin
		case state_reg is 
			when s0 => 
				P  <= 0;
				CC <= 0;
				CS <= 1;
				EN <= 1;
				LP <= 0;
			when s1 => 
				CC <= 1;
				CS <= 1;
				EN <= 1;			
			when s2 => 
				LP <= 1; 
			when s3 => 
				LP <= 0;
				EN <= 1;
				P <= not clk;
		end case;
	end process;

end architecture clocked_fsm_arch;