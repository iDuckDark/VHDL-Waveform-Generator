library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity triangle_entity is
    port ( 
        address : in std_logic_vector(6 downto 0);
        data : out real 
    );
end entity triangle_entity;

architecture triangle_arch of triangle_entity is
    type mem is array ( 0 to 99) of real;
    constant my_rom : mem := (
        0 =>-1.0,
        1 =>-0.980000000000000,
        2 =>-0.960000000000000,
        3 =>-0.940000000000000,
        4 =>-0.920000000000000,
        5 =>-0.900000000000000,
        6 =>-0.880000000000000,
        7 =>-0.860000000000000,
        8 =>-0.840000000000000,
        9 =>-0.820000000000000,
        10 =>-0.800000000000000,
        11 =>-0.780000000000000,
        12 =>-0.760000000000000,
        13 =>-0.740000000000000,
        14 =>-0.720000000000000,
        15 =>-0.700000000000000,
        16 =>-0.680000000000000,
        17 =>-0.660000000000000,
        18 =>-0.640000000000000,
        19 =>-0.620000000000000,
        20 =>-0.600000000000000,
        21 =>-0.580000000000000,
        22 =>-0.560000000000000,
        23 =>-0.540000000000000,
        24 =>-0.520000000000000,
        25 =>-0.500000000000000,
        26 =>-0.480000000000000,
        27 =>-0.460000000000000,
        28 =>-0.440000000000000,
        29 =>-0.420000000000000,
        30 =>-0.400000000000000,
        31 =>-0.380000000000000,
        32 =>-0.360000000000000,
        33 =>-0.340000000000000,
        34 =>-0.320000000000000,
        35 =>-0.300000000000000,
        36 =>-0.280000000000000,
        37 =>-0.260000000000000,
        38 =>-0.240000000000000,
        39 =>-0.220000000000000,
        40 =>-0.200000000000000,
        41 =>-0.180000000000000,
        42 =>-0.160000000000000,
        43 =>-0.140000000000000,
        44 =>-0.120000000000000,
        45 =>-0.100000000000000,
        46 =>-0.0800000000000000,
        47 =>-0.0599999999999999,
        48 =>-0.0399999999999999,
        49 =>-0.0199999999999999,
        50 =>-2.22044604925031e-16,
        51 =>0.0199999999999998,
        52 =>0.0399999999999998,
        53 =>0.0600000000000001,
        54 =>0.0799999999999996,
        55 =>0.0999999999999996,
        56 =>0.120000000000000,
        57 =>0.140000000000000,
        58 =>0.160000000000000,
        59 =>0.180000000000000,
        60 =>0.200000000000000,
        61 =>0.220000000000000,
        62 =>0.240000000000000,
        63 =>0.260000000000000,
        64 =>0.280000000000000,
        65 =>0.300000000000000,
        66 =>0.320000000000000,
        67 =>0.340000000000000,
        68 =>0.360000000000000,
        69 =>0.380000000000000,
        70 =>0.400000000000000,
        71 =>0.420000000000000,
        72 =>0.440000000000000,
        73 =>0.460000000000000,
        74 =>0.480000000000000,
        75 =>0.500000000000000,
        76 =>0.520000000000000,
        77 =>0.540000000000000,
        78 =>0.560000000000000,
        79 =>0.580000000000000,
        80 =>0.600000000000000,
        81 =>0.620000000000000,
        82 =>0.640000000000000,
        83 =>0.660000000000000,
        84 =>0.680000000000000,
        85 =>0.700000000000000,
        86 =>0.720000000000000,
        87 =>0.740000000000000,
        88 =>0.760000000000000,
        89 =>0.780000000000000,
        90 =>0.800000000000000,
        91 =>0.820000000000000,
        92 =>0.840000000000000,
        93 =>0.860000000000000,
        94 =>0.880000000000000,
        95 =>0.900000000000000,
        96 =>0.920000000000000,
        97 =>0.940000000000000,
        98 =>0.960000000000000,
        99 =>0.980000000000000);

    begin
        process (address)
        begin
          case address is
            when "0000000" => data <= my_rom(0);
            when "0000001" => data <= my_rom(1);
            when "0000010" => data <= my_rom(2);
            when "0000011" => data <= my_rom(3);
            when "0000100" => data <= my_rom(4);
            when "0000101" => data <= my_rom(5);
            when "0000110" => data <= my_rom(6);
            when "0000111" => data <= my_rom(7);
            when "0001000" => data <= my_rom(8);
            when "0001001" => data <= my_rom(9);
            when "0001010" => data <= my_rom(10);
            when "0001011" => data <= my_rom(11);
            when "0001100" => data <= my_rom(12);
            when "0001101" => data <= my_rom(13);
            when "0001110" => data <= my_rom(14);
            when "0001111" => data <= my_rom(15);
            when "0010000" => data <= my_rom(16);
            when "0010001" => data <= my_rom(17);
            when "0010010" => data <= my_rom(18);
            when "0010011" => data <= my_rom(19);
            when "0010100" => data <= my_rom(20);
            when "0010101" => data <= my_rom(21);
            when "0010110" => data <= my_rom(22);
            when "0010111" => data <= my_rom(23);
            when "0011000" => data <= my_rom(24);
            when "0011001" => data <= my_rom(25);
            when "0011010" => data <= my_rom(26);
            when "0011011" => data <= my_rom(27);
            when "0011100" => data <= my_rom(28);
            when "0011101" => data <= my_rom(29);
            when "0011110" => data <= my_rom(30);
            when "0011111" => data <= my_rom(31);
            when "0100000" => data <= my_rom(32);
            when "0100001" => data <= my_rom(33);
            when "0100010" => data <= my_rom(34);
            when "0100011" => data <= my_rom(35);
            when "0100100" => data <= my_rom(36);
            when "0100101" => data <= my_rom(37);
            when "0100110" => data <= my_rom(38);
            when "0100111" => data <= my_rom(39);
            when "0101000" => data <= my_rom(40);
            when "0101001" => data <= my_rom(41);
            when "0101010" => data <= my_rom(42);
            when "0101011" => data <= my_rom(43);
            when "0101100" => data <= my_rom(44);
            when "0101101" => data <= my_rom(45);
            when "0101110" => data <= my_rom(46);
            when "0101111" => data <= my_rom(47);
            when "0110000" => data <= my_rom(48);
            when "0110001" => data <= my_rom(49);
            when "0110010" => data <= my_rom(50);
            when "0110011" => data <= my_rom(51);
            when "0110100" => data <= my_rom(52);
            when "0110101" => data <= my_rom(53);
            when "0110110" => data <= my_rom(54);
            when "0110111" => data <= my_rom(55);
            when "0111000" => data <= my_rom(56);
            when "0111001" => data <= my_rom(57);
            when "0111010" => data <= my_rom(58);
            when "0111011" => data <= my_rom(59);
            when "0111100" => data <= my_rom(60);
            when "0111101" => data <= my_rom(61);
            when "0111110" => data <= my_rom(62);
            when "0111111" => data <= my_rom(63);
            when "1000000" => data <= my_rom(64);
            when "1000001" => data <= my_rom(65);
            when "1000010" => data <= my_rom(66);
            when "1000011" => data <= my_rom(67);
            when "1000100" => data <= my_rom(68);
            when "1000101" => data <= my_rom(69);
            when "1000110" => data <= my_rom(70);
            when "1000111" => data <= my_rom(71);
            when "1001000" => data <= my_rom(72);
            when "1001001" => data <= my_rom(73);
            when "1001010" => data <= my_rom(74);
            when "1001011" => data <= my_rom(75);
            when "1001100" => data <= my_rom(76);
            when "1001101" => data <= my_rom(77);
            when "1001110" => data <= my_rom(78);
            when "1001111" => data <= my_rom(79);
            when "1010000" => data <= my_rom(80);
            when "1010001" => data <= my_rom(81);
            when "1010010" => data <= my_rom(82);
            when "1010011" => data <= my_rom(83);
            when "1010100" => data <= my_rom(84);
            when "1010101" => data <= my_rom(85);
            when "1010110" => data <= my_rom(86);
            when "1010111" => data <= my_rom(87);
            when "1011000" => data <= my_rom(88);
            when "1011001" => data <= my_rom(89);
            when "1011010" => data <= my_rom(90);
            when "1011011" => data <= my_rom(91);
            when "1011100" => data <= my_rom(92);
            when "1011101" => data <= my_rom(93);
            when "1011110" => data <= my_rom(94);
            when "1011111" => data <= my_rom(95);
            when "1100000" => data <= my_rom(96);
            when "1100001" => data <= my_rom(97);
            when "1100010" => data <= my_rom(98);
            when "1100011" => data <= my_rom(99);
            when others => data <= 0.0;
          end case;
      end process;
end triangle_arch;
        