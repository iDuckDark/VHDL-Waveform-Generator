
    library ieee;
    use ieee.std_logic_1164.all;

    entity cos is
      port ( address : in std_logic_vector(6 downto 0);
             data : out real );
    end entity cos;

    architecture cos_arch of cos is
      type mem is array ( 0 to 99) of real;
      constant my_rom : mem := (
       0 =>1.0,
 1 =>0.998026728428272,
 2 =>0.992114701314478,
 3 =>0.982287250728689,
 4 =>0.968583161128631,
 5 =>0.951056516295154,
 6 =>0.929776485888251,
 7 =>0.904827052466020,
 8 =>0.876306680043864,
 9 =>0.844327925502015,
 10 =>0.809016994374948,
 11 =>0.770513242775789,
 12 =>0.728968627421412,
 13 =>0.684547105928689,
 14 =>0.637423989748690,
 15 =>0.587785252292473,
 16 =>0.535826794978997,
 17 =>0.481753674101715,
 18 =>0.425779291565073,
 19 =>0.368124552684678,
 20 =>0.309016994374947,
 21 =>0.248689887164855,
 22 =>0.187381314585725,
 23 =>0.125333233564304,
 24 =>0.0627905195293133,
 25 =>6.12323399573677e-17,
 26 =>-0.0627905195293134,
 27 =>-0.125333233564304,
 28 =>-0.187381314585725,
 29 =>-0.248689887164855,
 30 =>-0.309016994374947,
 31 =>-0.368124552684678,
 32 =>-0.425779291565073,
 33 =>-0.481753674101715,
 34 =>-0.535826794978996,
 35 =>-0.587785252292473,
 36 =>-0.637423989748690,
 37 =>-0.684547105928689,
 38 =>-0.728968627421411,
 39 =>-0.770513242775789,
 40 =>-0.809016994374947,
 41 =>-0.844327925502015,
 42 =>-0.876306680043864,
 43 =>-0.904827052466020,
 44 =>-0.929776485888251,
 45 =>-0.951056516295154,
 46 =>-0.968583161128631,
 47 =>-0.982287250728689,
 48 =>-0.992114701314478,
 49 =>-0.998026728428272,
 50 =>-1.0,
 51 =>-0.998026728428272,
 52 =>-0.992114701314478,
 53 =>-0.982287250728689,
 54 =>-0.968583161128631,
 55 =>-0.951056516295154,
 56 =>-0.929776485888252,
 57 =>-0.904827052466020,
 58 =>-0.876306680043864,
 59 =>-0.844327925502015,
 60 =>-0.809016994374948,
 61 =>-0.770513242775790,
 62 =>-0.728968627421412,
 63 =>-0.684547105928689,
 64 =>-0.637423989748690,
 65 =>-0.587785252292474,
 66 =>-0.535826794978997,
 67 =>-0.481753674101715,
 68 =>-0.425779291565073,
 69 =>-0.368124552684679,
 70 =>-0.309016994374948,
 71 =>-0.248689887164856,
 72 =>-0.187381314585726,
 73 =>-0.125333233564305,
 74 =>-0.0627905195293141,
 75 =>-1.83697019872103e-16,
 76 =>0.0627905195293128,
 77 =>0.125333233564303,
 78 =>0.187381314585724,
 79 =>0.248689887164854,
 80 =>0.309016994374946,
 81 =>0.368124552684677,
 82 =>0.425779291565072,
 83 =>0.481753674101715,
 84 =>0.535826794978996,
 85 =>0.587785252292472,
 86 =>0.637423989748689,
 87 =>0.684547105928688,
 88 =>0.728968627421411,
 89 =>0.770513242775789,
 90 =>0.809016994374947,
 91 =>0.844327925502015,
 92 =>0.876306680043864,
 93 =>0.904827052466019,
 94 =>0.929776485888251,
 95 =>0.951056516295154,
 96 =>0.968583161128631,
 97 =>0.982287250728689,
 98 =>0.992114701314478,
 99 =>0.998026728428272);

    begin
       process (address)
       begin
         case address is
         when "0000000" => data <= my_rom(0);
when "0000001" => data <= my_rom(1);
when "0000010" => data <= my_rom(2);
when "0000011" => data <= my_rom(3);
when "0000100" => data <= my_rom(4);
when "0000101" => data <= my_rom(5);
when "0000110" => data <= my_rom(6);
when "0000111" => data <= my_rom(7);
when "0001000" => data <= my_rom(8);
when "0001001" => data <= my_rom(9);
when "0001010" => data <= my_rom(10);
when "0001011" => data <= my_rom(11);
when "0001100" => data <= my_rom(12);
when "0001101" => data <= my_rom(13);
when "0001110" => data <= my_rom(14);
when "0001111" => data <= my_rom(15);
when "0010000" => data <= my_rom(16);
when "0010001" => data <= my_rom(17);
when "0010010" => data <= my_rom(18);
when "0010011" => data <= my_rom(19);
when "0010100" => data <= my_rom(20);
when "0010101" => data <= my_rom(21);
when "0010110" => data <= my_rom(22);
when "0010111" => data <= my_rom(23);
when "0011000" => data <= my_rom(24);
when "0011001" => data <= my_rom(25);
when "0011010" => data <= my_rom(26);
when "0011011" => data <= my_rom(27);
when "0011100" => data <= my_rom(28);
when "0011101" => data <= my_rom(29);
when "0011110" => data <= my_rom(30);
when "0011111" => data <= my_rom(31);
when "0100000" => data <= my_rom(32);
when "0100001" => data <= my_rom(33);
when "0100010" => data <= my_rom(34);
when "0100011" => data <= my_rom(35);
when "0100100" => data <= my_rom(36);
when "0100101" => data <= my_rom(37);
when "0100110" => data <= my_rom(38);
when "0100111" => data <= my_rom(39);
when "0101000" => data <= my_rom(40);
when "0101001" => data <= my_rom(41);
when "0101010" => data <= my_rom(42);
when "0101011" => data <= my_rom(43);
when "0101100" => data <= my_rom(44);
when "0101101" => data <= my_rom(45);
when "0101110" => data <= my_rom(46);
when "0101111" => data <= my_rom(47);
when "0110000" => data <= my_rom(48);
when "0110001" => data <= my_rom(49);
when "0110010" => data <= my_rom(50);
when "0110011" => data <= my_rom(51);
when "0110100" => data <= my_rom(52);
when "0110101" => data <= my_rom(53);
when "0110110" => data <= my_rom(54);
when "0110111" => data <= my_rom(55);
when "0111000" => data <= my_rom(56);
when "0111001" => data <= my_rom(57);
when "0111010" => data <= my_rom(58);
when "0111011" => data <= my_rom(59);
when "0111100" => data <= my_rom(60);
when "0111101" => data <= my_rom(61);
when "0111110" => data <= my_rom(62);
when "0111111" => data <= my_rom(63);
when "1000000" => data <= my_rom(64);
when "1000001" => data <= my_rom(65);
when "1000010" => data <= my_rom(66);
when "1000011" => data <= my_rom(67);
when "1000100" => data <= my_rom(68);
when "1000101" => data <= my_rom(69);
when "1000110" => data <= my_rom(70);
when "1000111" => data <= my_rom(71);
when "1001000" => data <= my_rom(72);
when "1001001" => data <= my_rom(73);
when "1001010" => data <= my_rom(74);
when "1001011" => data <= my_rom(75);
when "1001100" => data <= my_rom(76);
when "1001101" => data <= my_rom(77);
when "1001110" => data <= my_rom(78);
when "1001111" => data <= my_rom(79);
when "1010000" => data <= my_rom(80);
when "1010001" => data <= my_rom(81);
when "1010010" => data <= my_rom(82);
when "1010011" => data <= my_rom(83);
when "1010100" => data <= my_rom(84);
when "1010101" => data <= my_rom(85);
when "1010110" => data <= my_rom(86);
when "1010111" => data <= my_rom(87);
when "1011000" => data <= my_rom(88);
when "1011001" => data <= my_rom(89);
when "1011010" => data <= my_rom(90);
when "1011011" => data <= my_rom(91);
when "1011100" => data <= my_rom(92);
when "1011101" => data <= my_rom(93);
when "1011110" => data <= my_rom(94);
when "1011111" => data <= my_rom(95);
when "1100000" => data <= my_rom(96);
when "1100001" => data <= my_rom(97);
when "1100010" => data <= my_rom(98);
when "1100011" => data <= my_rom(99);

               when others => data <= 0.0;
                 end case;
          end process;
        end cos_arch;
        